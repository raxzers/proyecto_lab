magic
tech scmos
timestamp 1684113152
<< nwell >>
rect -16 -5 30 24
<< polysilicon >>
rect -4 9 0 26
rect 12 9 16 26
rect -4 -22 0 2
rect 12 -22 16 2
rect -4 -30 0 -28
rect 12 -30 16 -28
<< ndiffusion >>
rect -8 -28 -4 -22
rect 0 -28 12 -22
rect 16 -28 20 -22
<< pdiffusion >>
rect -8 2 -4 9
rect 0 2 4 9
rect 8 2 12 9
rect 16 2 20 9
<< metal1 >>
rect -4 30 0 37
rect 12 30 16 37
rect -12 18 -11 23
rect -6 18 4 23
rect 8 18 18 23
rect 23 18 38 23
rect -12 -6 -8 9
rect 4 2 8 18
rect 20 -6 24 9
rect -12 -11 37 -6
rect 20 -22 24 -11
rect -12 -35 -8 -28
rect -12 -39 -7 -35
rect -3 -39 3 -35
rect 7 -39 12 -35
rect 16 -39 24 -35
<< ntransistor >>
rect -4 -28 0 -22
rect 12 -28 16 -22
<< ptransistor >>
rect -4 2 0 9
rect 12 2 16 9
<< polycontact >>
rect -4 26 0 30
rect 12 26 16 30
<< ndcontact >>
rect -12 -28 -8 -22
rect 20 -28 24 -22
<< pdcontact >>
rect -12 2 -8 9
rect 4 2 8 9
rect 20 2 24 9
<< psubstratepcontact >>
rect -7 -39 -3 -35
rect 3 -39 7 -35
rect 12 -39 16 -35
<< nsubstratencontact >>
rect -11 18 -6 23
rect 4 18 8 23
rect 18 18 23 23
<< labels >>
rlabel metal1 -4 37 0 37 5 In1
rlabel metal1 12 37 16 37 5 In2
rlabel metal1 37 -11 37 -6 7 out
rlabel metal1 23 -37 23 -37 1 gnd!
rlabel metal1 35 21 35 21 7 vdd!
<< end >>
