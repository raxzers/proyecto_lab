magic
tech scmos
timestamp 1683997466
<< nwell >>
rect 3 0 33 26
<< polysilicon >>
rect 15 14 17 16
rect 15 -10 17 6
rect 15 -16 17 -14
<< ndiffusion >>
rect 14 -14 15 -10
rect 17 -14 18 -10
<< pdiffusion >>
rect 14 6 15 14
rect 17 6 18 14
<< metal1 >>
rect 3 18 7 22
rect 11 18 15 22
rect 19 18 23 22
rect 27 18 33 22
rect 10 14 14 18
rect 18 -3 22 6
rect 3 -7 11 -3
rect 18 -7 33 -3
rect 18 -10 22 -7
rect 10 -18 14 -14
rect 3 -22 7 -18
rect 11 -22 15 -18
rect 19 -22 23 -18
rect 27 -22 33 -18
<< ntransistor >>
rect 15 -14 17 -10
<< ptransistor >>
rect 15 6 17 14
<< polycontact >>
rect 11 -7 15 -3
<< ndcontact >>
rect 10 -14 14 -10
rect 18 -14 22 -10
<< pdcontact >>
rect 10 6 14 14
rect 18 6 22 14
<< psubstratepcontact >>
rect 7 -22 11 -18
rect 15 -22 19 -18
rect 23 -22 27 -18
<< nsubstratencontact >>
rect 7 18 11 22
rect 15 18 19 22
rect 23 18 27 22
<< labels >>
rlabel metal1 31 20 31 20 7 vdd!
rlabel metal1 30 -20 30 -20 8 gnd!
rlabel metal1 3 -7 3 -3 3 in
rlabel metal1 33 -7 33 -3 7 out
<< end >>
